`timescale 1ns / 1ps

module DUT
    (
        input Enable,
        input Reset,
        input Data,
        output Q
    );

     wire Q1;
     
     
     
     endmodule